module ledtest(output logic s);

	assign s = 1;
endmodule